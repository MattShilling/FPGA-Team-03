// unfinished
module IR_decoder(
input logic [15:0] dec;
input logic clk; 
);

endmodule
